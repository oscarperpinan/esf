*Celula

.subckt celula 303 300 302 310 

*Entre 300 y 301 está la fuente de corriente (de 300 a 301), 
*Fuente de corriente dependiente de la radiación (fuente de tensión)
*Entre 302(+) y 310(-) se aplica la entrada de radiación
*La salida se produce entre 303(+) y 300 (-)
*Isc depende de la radiación, que estará en kW/m2 (1 kW/m2 equivale a Isc)

grad 300 301 302 310 dc 4.3

d1 301 300 diode1
.model diode1 d is=1e-6 n=1.5

Rsh 301 300 {rsh}
Rs 301 303 {rs}

.ends

xcelD 6 5 102 100 celula rs=1e-4 rsh=1000
xcel5 5 4 101 100 celula rs=1e-4 rsh=1000
xcel4 4 3 101 100 celula rs=1e-4 rsh=1000
xcel3 3 2 101 100 celula rs=1e-4 rsh=1000
xcel2 2 1 101 100 celula rs=1e-4 rsh=1000
xcel1 1 0 101 100 celula rs=1e-4 rsh=1000

vbias 6 0 dc 0
vrad1 101 100 dc 1
vrad2 102 100 dc 0.99

*.print dc r(Rs.xcelD) v(6) v(5) v(1) i(Rs.xcelD)
*.dc Rsh.xcelD 1 10000 decade 3 Rs.xcelD 1e-4 1e-2 decade 1 vbias 0 1.2 0.01 >DispersionResistencias.dat
.print dc i(Rsh.xcelD) i(Rsh.xcel1) v(vbias) i(vbias) v(5) v(1) 
.dc Rsh.xcelD 1 10000 decade 3 vbias 0 3.6 0.01 >DispersionResistencias.dat



.end
