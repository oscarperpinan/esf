*Estudio de la influencia de la resistencia serie y resitencia paralelo en la
*característica I-V de una céula solar

.subckt celula 303 300 302 310 
.param rs=1 rsh=1

*Entre 300 y 301 está la fuente de corriente (de 300 a 301), 
*Fuente de corriente dependiente de la radiación (fuente de tensión)
*Entre 302(+) y 310(-) se aplica la entrada de radiación
*La salida se produce entre 303(+) y 300 (-)
*Isc depende de la radiación, que estará en kW/m2 (1 kW/m2 equivale a Isc)

grad 300 301 302 310 dc 4.3

d1 301 300 diode1
.model diode1 d is=1e-6 n=1.5

Rsh 301 300 {rsh}
Rs 301 303 {rs}

.ends

xcel1 1 0 101 100 celula rs=1e-4 rsh=100

vbias 1 0 dc 0
vrad1 101 100 dc 1

.print dc v(1) i(Rs.xcel1)
.dc Rs.xcel1 1e-4 1e-2 decade 1 vbias 0 0.6 0.01 >InfluenciaResistenciaSerie.dat
.dc Rsh.xcel1 1 100 decade 1 vbias 0 0.6 0.01 >InfluenciaResistenciaParalelo.dat



.end
