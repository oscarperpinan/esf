.subckt cell_2 300 303 302 
.param area=1 j0=1 jsc=1 j02=1 rs=1 rsh=1

girrad 301 300 302 300 value={(jsc/1000)*v(302)*area}

d1 301 300 diode
.model diode d(is={j0*area})

d2 301 300 diode2
.model diode2 d(is={j02*area}, n=2)

Rs 301 300 {rs}
Rsh 301 302 {rsh}

.ends

xcell2 0 31 32 cell_2 
*.param area=126.6 j0=1e11 j02=1E-9 jsc=0.0343 rs={RS} rsh=100000
*.param RS=1
vbias 31 0 dc 0
virrad 32 0 dc 1000

.print dc i(vbias)
.dc vbias 0.1 0.6 0.01 >cell_2.dat
*.step param RS list 0.0001 0.001 0.01 0.1 1
*.probe

.end